// mux4x1.v, 4x1 muxer, gate synthesis
//
// how to compile: ~changw/ivl/bin/iverilog decoder1x2.v
// how to run: ./a.out

module MuxMod(s1, s0, d0, d1, d2, d3, o); // module definition
   input s1, s0, d0, d1, d2, d3;
   output o;

   wire s1_inv, s0_inv, and0, and1, and2, and3;

   not(s1_inv, s1);
   not(s0_inv, s0);

   and(and0, d0, s0_inv, s1_inv);
   and(and1, d1, s0, s1_inv);
   and(and2, d2, s0_inv, s1);
   and(and3, d3, s0, s1);
   or(o, and0, and1, and2, and3);

endmodule

module TestMod; 
   reg s1, s0, d0, d1, d2, d3;       
   wire o;                          

   MuxMod my_muxer(s1, s0, d0, d1, d2, d3, o); // create instance

   initial begin
      $monitor("%0d\t%b\t%b\t%b\t%b\t%b\t%b\t%b", $time, s1, s0, d0, d1, d2, d3, o);
      $display("Time\ts1\ts0\td0\td1\td1\td1\to");
      $display("-----------------------------------------------------------------");
   end

   initial begin
      s1 = 0; s0 = 0; d0 = 0; d1 = 0; d2 = 0; d3 = 0;
      #1;
      s1 = 0; s0 = 0; d0 = 0; d1 = 0; d2 = 0; d3 = 1;
      #1;
      s1 = 0; s0 = 0; d0 = 0; d1 = 0; d2 = 1; d3 = 0;
      #1;
      s1 = 0; s0 = 0; d0 = 0; d1 = 0; d2 = 1; d3 = 1;
      #1;
      s1 = 0; s0 = 0; d0 = 0; d1 = 1; d2 = 0; d3 = 0;
      #1;
      s1 = 0; s0 = 0; d0 = 0; d1 = 1; d2 = 0; d3 = 1;
      #1;
      s1 = 0; s0 = 0; d0 = 0; d1 = 1; d2 = 1; d3 = 0;
      #1;
      s1 = 0; s0 = 0; d0 = 0; d1 = 1; d2 = 1; d3 = 1;
      #1;
      s1 = 0; s0 = 0; d0 = 1; d1 = 0; d2 = 0; d3 = 0;
      #1;
      s1 = 0; s0 = 0; d0 = 1; d1 = 0; d2 = 0; d3 = 1;
      #1;
      s1 = 0; s0 = 0; d0 = 1; d1 = 0; d2 = 1; d3 = 0;
      #1;
      s1 = 0; s0 = 0; d0 = 1; d1 = 0; d2 = 1; d3 = 1;
      #1;
      s1 = 0; s0 = 0; d0 = 1; d1 = 1; d2 = 0; d3 = 0;
      #1;
      s1 = 0; s0 = 0; d0 = 1; d1 = 1; d2 = 0; d3 = 1;
      #1;
      s1 = 0; s0 = 0; d0 = 1; d1 = 1; d2 = 1; d3 = 0;
      #1;
      s1 = 0; s0 = 0; d0 = 1; d1 = 1; d2 = 1; d3 = 1;
      #1;
      s1 = 0; s0 = 1; d0 = 0; d1 = 0; d2 = 0; d3 = 0;
      #1;
      s1 = 0; s0 = 1; d0 = 0; d1 = 0; d2 = 0; d3 = 1;
      #1;
      s1 = 0; s0 = 1; d0 = 0; d1 = 0; d2 = 1; d3 = 0;
      #1;
      s1 = 0; s0 = 1; d0 = 0; d1 = 0; d2 = 1; d3 = 1;
      #1;
      s1 = 0; s0 = 1; d0 = 0; d1 = 1; d2 = 0; d3 = 0;
      #1;
      s1 = 0; s0 = 1; d0 = 0; d1 = 1; d2 = 0; d3 = 1;
      #1;
      s1 = 0; s0 = 1; d0 = 0; d1 = 1; d2 = 1; d3 = 0;
      #1;
      s1 = 0; s0 = 1; d0 = 0; d1 = 1; d2 = 1; d3 = 1;
      #1;
      s1 = 0; s0 = 1; d0 = 1; d1 = 0; d2 = 0; d3 = 0;
      #1;
      s1 = 0; s0 = 1; d0 = 1; d1 = 0; d2 = 0; d3 = 1;
      #1;
      s1 = 0; s0 = 1; d0 = 1; d1 = 0; d2 = 1; d3 = 0;
      #1;
      s1 = 0; s0 = 1; d0 = 1; d1 = 0; d2 = 1; d3 = 1;
      #1;
      s1 = 0; s0 = 1; d0 = 1; d1 = 1; d2 = 0; d3 = 0;
      #1;
      s1 = 0; s0 = 1; d0 = 1; d1 = 1; d2 = 0; d3 = 1;
      #1;
      s1 = 0; s0 = 1; d0 = 1; d1 = 1; d2 = 1; d3 = 0;
      #1;
      s1 = 0; s0 = 1; d0 = 1; d1 = 1; d2 = 1; d3 = 1;
      #1;
      s1 = 1; s0 = 0; d0 = 0; d1 = 0; d2 = 0; d3 = 0;
      #1;
      s1 = 1; s0 = 0; d0 = 0; d1 = 0; d2 = 0; d3 = 1;
      #1;
      s1 = 1; s0 = 0; d0 = 0; d1 = 0; d2 = 1; d3 = 0;
      #1;
      s1 = 1; s0 = 0; d0 = 0; d1 = 0; d2 = 1; d3 = 1;
      #1;
      s1 = 1; s0 = 0; d0 = 0; d1 = 1; d2 = 0; d3 = 0;
      #1;
      s1 = 1; s0 = 0; d0 = 0; d1 = 1; d2 = 0; d3 = 1;
      #1;
      s1 = 1; s0 = 0; d0 = 0; d1 = 1; d2 = 1; d3 = 0;
      #1;
      s1 = 1; s0 = 0; d0 = 0; d1 = 1; d2 = 1; d3 = 1;
      #1;
      s1 = 1; s0 = 0; d0 = 1; d1 = 0; d2 = 0; d3 = 0;
      #1;
      s1 = 1; s0 = 0; d0 = 1; d1 = 0; d2 = 0; d3 = 1;
      #1;
      s1 = 1; s0 = 0; d0 = 1; d1 = 0; d2 = 1; d3 = 0;
      #1;
      s1 = 1; s0 = 0; d0 = 1; d1 = 0; d2 = 1; d3 = 1;
      #1;
      s1 = 1; s0 = 0; d0 = 1; d1 = 1; d2 = 0; d3 = 0;
      #1;
      s1 = 1; s0 = 0; d0 = 1; d1 = 1; d2 = 0; d3 = 1;
      #1;
      s1 = 1; s0 = 0; d0 = 1; d1 = 1; d2 = 1; d3 = 0;
      #1;
      s1 = 1; s0 = 0; d0 = 1; d1 = 1; d2 = 1; d3 = 1;
      #1;
      s1 = 1; s0 = 1; d0 = 0; d1 = 0; d2 = 0; d3 = 0;
      #1;
      s1 = 1; s0 = 1; d0 = 0; d1 = 0; d2 = 0; d3 = 1;
      #1;
      s1 = 1; s0 = 1; d0 = 0; d1 = 0; d2 = 1; d3 = 0;
      #1;
      s1 = 1; s0 = 1; d0 = 0; d1 = 0; d2 = 1; d3 = 1;
      #1;
      s1 = 1; s0 = 1; d0 = 0; d1 = 1; d2 = 0; d3 = 0;
      #1;
      s1 = 1; s0 = 1; d0 = 0; d1 = 1; d2 = 0; d3 = 1;
      #1;
      s1 = 1; s0 = 1; d0 = 0; d1 = 1; d2 = 1; d3 = 0;
      #1;
      s1 = 1; s0 = 1; d0 = 0; d1 = 1; d2 = 1; d3 = 1;
      #1;
      s1 = 1; s0 = 1; d0 = 1; d1 = 0; d2 = 0; d3 = 0;
      #1;
      s1 = 1; s0 = 1; d0 = 1; d1 = 0; d2 = 0; d3 = 1;
      #1;
      s1 = 1; s0 = 1; d0 = 1; d1 = 0; d2 = 1; d3 = 0;
      #1;
      s1 = 1; s0 = 1; d0 = 1; d1 = 0; d2 = 1; d3 = 1;
      #1;
      s1 = 1; s0 = 1; d0 = 1; d1 = 1; d2 = 0; d3 = 0;
      #1;
      s1 = 1; s0 = 1; d0 = 1; d1 = 1; d2 = 0; d3 = 1;
      #1;
      s1 = 1; s0 = 1; d0 = 1; d1 = 1; d2 = 1; d3 = 0;
      #1;
      s1 = 1; s0 = 1; d0 = 1; d1 = 1; d2 = 1; d3 = 1;      
      #1;
   end
endmodule
