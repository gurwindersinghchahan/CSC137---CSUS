// Edward Prokopik

module MuxMod( s, d, o);
    input [1:0] s;
    input [0:3] d;
    output o;

    wire [0:1] s_inv;
    wire [0:3] ands;

    not(s_inv[1], s[1]);
    not(s_inv[0], s[0]);
    and(ands[0], d[0], s_inv[1], s_inv[0]);
    and(ands[1], d[1], s_inv[1], s[0]);
    and(ands[2], d[2], s[1], s_inv[0]);
    and(ands[3], d[3], s[1], s[0]);
    or(o, ands[0], ands[1], ands[2], ands[3]);

endmodule

module TestMod;

   reg [0:1] s;
   reg [0:3] d;       
   wire o;                          

   MuxMod mux_n_mod (s, d, o); 

   initial begin
      $monitor("%0d\t%b\t%b\t%b",
             $time, s, d, o);
      $display("Time\ts\td\to");
      $display("-----------------------------------------------------------------");
   end

   initial begin
      s = 2'b00; d = 4'b0000; #1;
      s = 2'b00; d = 4'b0001; #1;
      s = 2'b00; d = 4'b0010; #1;
      s = 2'b00; d = 4'b0011; #1;
      s = 2'b00; d = 4'b0100; #1;
      s = 2'b00; d = 4'b0101; #1;
      s = 2'b00; d = 4'b0110; #1;
      s = 2'b00; d = 4'b0111; #1;
      s = 2'b00; d = 4'b1000; #1;
      s = 2'b00; d = 4'b1001; #1;
      s = 2'b00; d = 4'b1010; #1;
      s = 2'b00; d = 4'b1011; #1;
      s = 2'b00; d = 4'b1100; #1;
      s = 2'b00; d = 4'b1101; #1;
      s = 2'b00; d = 4'b1110; #1;
      s = 2'b00; d = 4'b1111; #1;

      s = 2'b01; d = 4'b0000; #1;
      s = 2'b01; d = 4'b0001; #1;
      s = 2'b01; d = 4'b0010; #1;
      s = 2'b01; d = 4'b0011; #1;
      s = 2'b01; d = 4'b0100; #1;
      s = 2'b01; d = 4'b0101; #1;
      s = 2'b01; d = 4'b0110; #1;
      s = 2'b01; d = 4'b0111; #1;
      s = 2'b01; d = 4'b1000; #1;
      s = 2'b01; d = 4'b1001; #1;
      s = 2'b01; d = 4'b1010; #1;
      s = 2'b01; d = 4'b1011; #1;
      s = 2'b01; d = 4'b1100; #1;
      s = 2'b01; d = 4'b1101; #1;
      s = 2'b01; d = 4'b1110; #1;
      s = 2'b01; d = 4'b1111; #1;

      s = 2'b10; d = 4'b0000; #1;
      s = 2'b10; d = 4'b0001; #1;
      s = 2'b10; d = 4'b0010; #1;
      s = 2'b10; d = 4'b0011; #1;
      s = 2'b10; d = 4'b0100; #1;
      s = 2'b10; d = 4'b0101; #1;
      s = 2'b10; d = 4'b0110; #1;
      s = 2'b10; d = 4'b0111; #1;
      s = 2'b10; d = 4'b1000; #1;
      s = 2'b10; d = 4'b1001; #1;
      s = 2'b10; d = 4'b1010; #1;
      s = 2'b10; d = 4'b1011; #1;
      s = 2'b10; d = 4'b1100; #1;
      s = 2'b10; d = 4'b1101; #1;
      s = 2'b10; d = 4'b1110; #1;
      s = 2'b10; d = 4'b1111; #1;

      s = 2'b11; d = 4'b0000; #1;
      s = 2'b11; d = 4'b0001; #1;
      s = 2'b11; d = 4'b0010; #1;
      s = 2'b11; d = 4'b0011; #1;
      s = 2'b11; d = 4'b0100; #1;
      s = 2'b11; d = 4'b0101; #1;
      s = 2'b11; d = 4'b0110; #1;
      s = 2'b11; d = 4'b0111; #1;
      s = 2'b11; d = 4'b1000; #1;
      s = 2'b11; d = 4'b1001; #1;
      s = 2'b11; d = 4'b1010; #1;
      s = 2'b11; d = 4'b1011; #1;
      s = 2'b11; d = 4'b1100; #1;
      s = 2'b11; d = 4'b1101; #1;
      s = 2'b11; d = 4'b1110; #1;
      s = 2'b11; d = 4'b1111; #1;

   end
endmodule